`timescale 1ns / 1ps

module ad9361_reg_test(clk,rst_n,index,cmd_datao );
    input clk;   
    input rst_n; 
    input[15:0] index;
    output[23:0] cmd_datao;
    reg[18:0] cmd_data;
    reg[23:0] cmd_datao;
    reg[18:0] waiting = {1'b1,10'hFFF,8'hFF};
    
    always @ (posedge clk)
        if(cmd_data == waiting)
            cmd_datao <= {1'b0,5'b11111,cmd_data[17:0]};
        else
            cmd_datao <= {cmd_data[18],5'b00000,cmd_data[17:0]};
    
    always @ (*) 
        begin
            case(index)
               -12'd2  :cmd_data={1'b1,10'hFFF,8'hFF};//set spi  --
               -12'd1  :cmd_data={1'b1,10'h000,8'h00};//set spi  --
                12'd0  :cmd_data={1'b1,10'h3DF,8'h01};
                12'd1  :cmd_data={1'b1,10'h2A6,8'h0E};
                12'd2  :cmd_data={1'b1,10'h2A8,8'h0E};
                12'd3  :cmd_data={1'b1,10'h2AB,8'h07};
                12'd4  :cmd_data={1'b1,10'h2AC,8'hFF};
                12'd5  :cmd_data={1'b1,10'h009,8'h17};
                12'd6  :cmd_data={1'b1,10'hFFF,8'hFF};
                12'd7  :cmd_data={1'b1,10'h045,8'h00};
                12'd8  :cmd_data={1'b1,10'h046,8'h06};
                12'd9  :cmd_data={1'b1,10'h048,8'hE8};
                12'd10  :cmd_data={1'b1,10'h049,8'h5B};
                12'd11  :cmd_data={1'b1,10'h04A,8'h35};
                12'd12  :cmd_data={1'b1,10'h04B,8'hE0};
                12'd13  :cmd_data={1'b1,10'h04E,8'h10};
                12'd14  :cmd_data={1'b1,10'h043,8'h00};
                12'd15  :cmd_data={1'b1,10'h042,8'h00};
                12'd16  :cmd_data={1'b1,10'h041,8'h00};
                12'd17  :cmd_data={1'b1,10'h044,8'h28};
                12'd18  :cmd_data={1'b1,10'h03F,8'h05};
                12'd19  :cmd_data={1'b1,10'h03F,8'h01};
                12'd20  :cmd_data={1'b1,10'h04C,8'h86};
                12'd21  :cmd_data={1'b1,10'h04D,8'h01};
                12'd22  :cmd_data={1'b1,10'h04D,8'h05};
                12'd23  :cmd_data={1'b0,10'h05E,8'h00};
                12'd24  :cmd_data={1'b1,10'h002,8'h04};
                12'd25  :cmd_data={1'b1,10'h003,8'h44};
                12'd26  :cmd_data={1'b1,10'h004,8'h03};
                12'd27  :cmd_data={1'b1,10'h00A,8'h02};
                12'd28  :cmd_data={1'b1,10'h010,8'hC8};
                12'd29  :cmd_data={1'b1,10'h011,8'h00};
                12'd30  :cmd_data={1'b1,10'h012,8'h10};
                12'd31  :cmd_data={1'b1,10'h006,8'h00};
                12'd32  :cmd_data={1'b1,10'h007,8'h00};
                12'd33  :cmd_data={1'b1,10'h03C,8'h23};
                12'd34  :cmd_data={1'b1,10'h03D,8'hFF};
                12'd35  :cmd_data={1'b1,10'h03E,8'h0F};
                12'd36  :cmd_data={1'b1,10'h018,8'h00};
                12'd37  :cmd_data={1'b1,10'h019,8'h00};
                12'd38  :cmd_data={1'b1,10'h01A,8'h00};
                12'd39  :cmd_data={1'b1,10'h01B,8'h00};
                12'd40  :cmd_data={1'b1,10'h023,8'hFF};
                12'd41  :cmd_data={1'b1,10'h026,8'h00};
                12'd42  :cmd_data={1'b1,10'h030,8'h00};
                12'd43  :cmd_data={1'b1,10'h031,8'h00};
                12'd44  :cmd_data={1'b1,10'h032,8'h00};
                12'd45  :cmd_data={1'b1,10'h033,8'h00};
                12'd46  :cmd_data={1'b1,10'h00B,8'h00};
                12'd47  :cmd_data={1'b1,10'h00C,8'h00};
                12'd48  :cmd_data={1'b1,10'h00D,8'h03};
                12'd49  :cmd_data={1'b1,10'h00F,8'h04};
                12'd50  :cmd_data={1'b1,10'h01C,8'h10};
                12'd51  :cmd_data={1'b1,10'h01D,8'h01};
                12'd52  :cmd_data={1'b1,10'h035,8'h00};
                12'd53  :cmd_data={1'b1,10'h036,8'hFF};
                12'd54  :cmd_data={1'b1,10'h03A,8'h13};
                12'd55  :cmd_data={1'b1,10'h020,8'h00};
                12'd56  :cmd_data={1'b1,10'h027,8'h03};
                12'd57  :cmd_data={1'b1,10'h028,8'h00};
                12'd58  :cmd_data={1'b1,10'h029,8'h00};
                12'd59  :cmd_data={1'b1,10'h02A,8'h00};
                12'd60  :cmd_data={1'b1,10'h02B,8'h00};
                12'd61  :cmd_data={1'b1,10'h02C,8'h00};
                12'd62  :cmd_data={1'b1,10'h02D,8'h00};
                12'd63  :cmd_data={1'b1,10'h02E,8'h00};
                12'd64  :cmd_data={1'b1,10'h02F,8'h00};
                12'd65  :cmd_data={1'b1,10'h261,8'h00};
                12'd66  :cmd_data={1'b1,10'h2A1,8'h00};
                12'd67  :cmd_data={1'b1,10'h248,8'h0B};
                12'd68  :cmd_data={1'b1,10'h288,8'h0B};
                12'd69  :cmd_data={1'b1,10'h246,8'h02};
                12'd70  :cmd_data={1'b1,10'h286,8'h02};
                12'd71  :cmd_data={1'b1,10'h249,8'h8E};
                12'd72  :cmd_data={1'b1,10'h289,8'h8E};
                12'd73  :cmd_data={1'b1,10'h23B,8'h80};
                12'd74  :cmd_data={1'b1,10'h27B,8'h80};
                12'd75  :cmd_data={1'b1,10'h243,8'h0D};
                12'd76  :cmd_data={1'b1,10'h283,8'h0D};
                12'd77  :cmd_data={1'b1,10'h23D,8'h00};
                12'd78  :cmd_data={1'b1,10'h27D,8'h00};
                12'd79  :cmd_data={1'b1,10'h015,8'h04};
                12'd80  :cmd_data={1'b1,10'h014,8'h05};
                12'd81  :cmd_data={1'b1,10'h013,8'h01};
                12'd82  :cmd_data={1'b0,10'h017,8'h00};
                12'd83  :cmd_data={1'b1,10'h23D,8'h04};
                12'd84  :cmd_data={1'b0,10'h244,8'h00};
                12'd85  :cmd_data={1'b1,10'h27D,8'h04};
                12'd86  :cmd_data={1'b0,10'h284,8'h00};
                12'd87  :cmd_data={1'b1,10'h23D,8'h00};
                12'd88  :cmd_data={1'b1,10'h27D,8'h00};
                12'd89  :cmd_data={1'b1,10'h23A,8'h4A};
                12'd90  :cmd_data={1'b1,10'h239,8'hC1};
                12'd91  :cmd_data={1'b1,10'h242,8'h17};
                12'd92  :cmd_data={1'b1,10'h238,8'h78};
                12'd93  :cmd_data={1'b1,10'h245,8'h00};
                12'd94  :cmd_data={1'b1,10'h251,8'h0E};
                12'd95  :cmd_data={1'b1,10'h250,8'h70};
                12'd96  :cmd_data={1'b1,10'h23B,8'h96};
                12'd97  :cmd_data={1'b1,10'h23E,8'hC3};
                12'd98  :cmd_data={1'b1,10'h23F,8'hEF};
                12'd99  :cmd_data={1'b1,10'h240,8'h0B};
                12'd100  :cmd_data={1'b1,10'h27A,8'h4A};
                12'd101  :cmd_data={1'b1,10'h279,8'hC1};
                12'd102  :cmd_data={1'b1,10'h282,8'h17};
                12'd103  :cmd_data={1'b1,10'h278,8'h78};
                12'd104  :cmd_data={1'b1,10'h285,8'h00};
                12'd105  :cmd_data={1'b1,10'h291,8'h0E};
                12'd106  :cmd_data={1'b1,10'h290,8'h70};
                12'd107  :cmd_data={1'b1,10'h27B,8'h96};
                12'd108  :cmd_data={1'b1,10'h27E,8'hC3};
                12'd109  :cmd_data={1'b1,10'h27F,8'hEF};
                12'd110  :cmd_data={1'b1,10'h280,8'h0B};
                12'd111  :cmd_data={1'b1,10'h233,8'hF5};
                12'd112  :cmd_data={1'b1,10'h234,8'hFF};
                12'd113  :cmd_data={1'b1,10'h235,8'h5F};
                12'd114  :cmd_data={1'b1,10'h232,8'h00};
                12'd115  :cmd_data={1'b1,10'h231,8'hB2};  // 3500 00AF 000000   3575 00B2 5FFFF5
                12'd116  :cmd_data={1'b1,10'h005,8'h00};
                12'd117  :cmd_data={1'b1,10'h273,8'hF5};
                12'd118  :cmd_data={1'b1,10'h274,8'hFF};
                12'd119  :cmd_data={1'b1,10'h275,8'h5F};
                12'd120  :cmd_data={1'b1,10'h272,8'h00};
                12'd121  :cmd_data={1'b1,10'h271,8'hB2};
                12'd122  :cmd_data={1'b1,10'h005,8'h00};
                12'd123  :cmd_data={1'b0,10'h247,8'h00};
                12'd124  :cmd_data={1'b0,10'h287,8'h00};
                12'd125  :cmd_data={1'b1,10'h13F,8'h02};
                12'd126  :cmd_data={1'b1,10'h138,8'h0F};
                12'd127  :cmd_data={1'b1,10'h139,8'h78};
                12'd128  :cmd_data={1'b1,10'h13A,8'h00};
                12'd129  :cmd_data={1'b1,10'h13B,8'h00};
                12'd130  :cmd_data={1'b1,10'h13F,8'h06};
                12'd131  :cmd_data={1'b1,10'h13C,8'h00};
                12'd132  :cmd_data={1'b1,10'h13C,8'h00};
                12'd133  :cmd_data={1'b1,10'h138,8'h0E};
                12'd134  :cmd_data={1'b1,10'h139,8'h74};
                12'd135  :cmd_data={1'b1,10'h13A,8'h00};
                12'd136  :cmd_data={1'b1,10'h13B,8'h0D};
                12'd137  :cmd_data={1'b1,10'h13F,8'h06};
                12'd138  :cmd_data={1'b1,10'h13C,8'h00};
                12'd139  :cmd_data={1'b1,10'h13C,8'h00};
                12'd140  :cmd_data={1'b1,10'h138,8'h0D};
                12'd141  :cmd_data={1'b1,10'h139,8'h70};
                12'd142  :cmd_data={1'b1,10'h13A,8'h00};
                12'd143  :cmd_data={1'b1,10'h13B,8'h15};
                12'd144  :cmd_data={1'b1,10'h13F,8'h06};
                12'd145  :cmd_data={1'b1,10'h13C,8'h00};
                12'd146  :cmd_data={1'b1,10'h13C,8'h00};
                12'd147  :cmd_data={1'b1,10'h138,8'h0C};
                12'd148  :cmd_data={1'b1,10'h139,8'h6C};
                12'd149  :cmd_data={1'b1,10'h13A,8'h00};
                12'd150  :cmd_data={1'b1,10'h13B,8'h1B};
                12'd151  :cmd_data={1'b1,10'h13F,8'h06};
                12'd152  :cmd_data={1'b1,10'h13C,8'h00};
                12'd153  :cmd_data={1'b1,10'h13C,8'h00};
                12'd154  :cmd_data={1'b1,10'h138,8'h0B};
                12'd155  :cmd_data={1'b1,10'h139,8'h68};
                12'd156  :cmd_data={1'b1,10'h13A,8'h00};
                12'd157  :cmd_data={1'b1,10'h13B,8'h21};
                12'd158  :cmd_data={1'b1,10'h13F,8'h06};
                12'd159  :cmd_data={1'b1,10'h13C,8'h00};
                12'd160  :cmd_data={1'b1,10'h13C,8'h00};
                12'd161  :cmd_data={1'b1,10'h138,8'h0A};
                12'd162  :cmd_data={1'b1,10'h139,8'h64};
                12'd163  :cmd_data={1'b1,10'h13A,8'h00};
                12'd164  :cmd_data={1'b1,10'h13B,8'h25};
                12'd165  :cmd_data={1'b1,10'h13F,8'h06};
                12'd166  :cmd_data={1'b1,10'h13C,8'h00};
                12'd167  :cmd_data={1'b1,10'h13C,8'h00};
                12'd168  :cmd_data={1'b1,10'h138,8'h09};
                12'd169  :cmd_data={1'b1,10'h139,8'h60};
                12'd170  :cmd_data={1'b1,10'h13A,8'h00};
                12'd171  :cmd_data={1'b1,10'h13B,8'h29};
                12'd172  :cmd_data={1'b1,10'h13F,8'h06};
                12'd173  :cmd_data={1'b1,10'h13C,8'h00};
                12'd174  :cmd_data={1'b1,10'h13C,8'h00};
                12'd175  :cmd_data={1'b1,10'h138,8'h08};
                12'd176  :cmd_data={1'b1,10'h139,8'h5C};
                12'd177  :cmd_data={1'b1,10'h13A,8'h00};
                12'd178  :cmd_data={1'b1,10'h13B,8'h2C};
                12'd179  :cmd_data={1'b1,10'h13F,8'h06};
                12'd180  :cmd_data={1'b1,10'h13C,8'h00};
                12'd181  :cmd_data={1'b1,10'h13C,8'h00};
                12'd182  :cmd_data={1'b1,10'h138,8'h07};
                12'd183  :cmd_data={1'b1,10'h139,8'h58};
                12'd184  :cmd_data={1'b1,10'h13A,8'h00};
                12'd185  :cmd_data={1'b1,10'h13B,8'h2F};
                12'd186  :cmd_data={1'b1,10'h13F,8'h06};
                12'd187  :cmd_data={1'b1,10'h13C,8'h00};
                12'd188  :cmd_data={1'b1,10'h13C,8'h00};
                12'd189  :cmd_data={1'b1,10'h138,8'h06};
                12'd190  :cmd_data={1'b1,10'h139,8'h54};
                12'd191  :cmd_data={1'b1,10'h13A,8'h00};
                12'd192  :cmd_data={1'b1,10'h13B,8'h31};
                12'd193  :cmd_data={1'b1,10'h13F,8'h06};
                12'd194  :cmd_data={1'b1,10'h13C,8'h00};
                12'd195  :cmd_data={1'b1,10'h13C,8'h00};
                12'd196  :cmd_data={1'b1,10'h138,8'h05};
                12'd197  :cmd_data={1'b1,10'h139,8'h50};
                12'd198  :cmd_data={1'b1,10'h13A,8'h00};
                12'd199  :cmd_data={1'b1,10'h13B,8'h33};
                12'd200  :cmd_data={1'b1,10'h13F,8'h06};
                12'd201  :cmd_data={1'b1,10'h13C,8'h00};
                12'd202  :cmd_data={1'b1,10'h13C,8'h00};
                12'd203  :cmd_data={1'b1,10'h138,8'h04};
                12'd204  :cmd_data={1'b1,10'h139,8'h4C};
                12'd205  :cmd_data={1'b1,10'h13A,8'h00};
                12'd206  :cmd_data={1'b1,10'h13B,8'h34};
                12'd207  :cmd_data={1'b1,10'h13F,8'h06};
                12'd208  :cmd_data={1'b1,10'h13C,8'h00};
                12'd209  :cmd_data={1'b1,10'h13C,8'h00};
                12'd210  :cmd_data={1'b1,10'h138,8'h03};
                12'd211  :cmd_data={1'b1,10'h139,8'h48};
                12'd212  :cmd_data={1'b1,10'h13A,8'h00};
                12'd213  :cmd_data={1'b1,10'h13B,8'h35};
                12'd214  :cmd_data={1'b1,10'h13F,8'h06};
                12'd215  :cmd_data={1'b1,10'h13C,8'h00};
                12'd216  :cmd_data={1'b1,10'h13C,8'h00};
                12'd217  :cmd_data={1'b1,10'h138,8'h02};
                12'd218  :cmd_data={1'b1,10'h139,8'h30};
                12'd219  :cmd_data={1'b1,10'h13A,8'h00};
                12'd220  :cmd_data={1'b1,10'h13B,8'h3A};
                12'd221  :cmd_data={1'b1,10'h13F,8'h06};
                12'd222  :cmd_data={1'b1,10'h13C,8'h00};
                12'd223  :cmd_data={1'b1,10'h13C,8'h00};
                12'd224  :cmd_data={1'b1,10'h138,8'h01};
                12'd225  :cmd_data={1'b1,10'h139,8'h18};
                12'd226  :cmd_data={1'b1,10'h13A,8'h00};
                12'd227  :cmd_data={1'b1,10'h13B,8'h3D};
                12'd228  :cmd_data={1'b1,10'h13F,8'h06};
                12'd229  :cmd_data={1'b1,10'h13C,8'h00};
                12'd230  :cmd_data={1'b1,10'h13C,8'h00};
                12'd231  :cmd_data={1'b1,10'h138,8'h00};
                12'd232  :cmd_data={1'b1,10'h139,8'h00};
                12'd233  :cmd_data={1'b1,10'h13A,8'h00};
                12'd234  :cmd_data={1'b1,10'h13B,8'h3E};
                12'd235  :cmd_data={1'b1,10'h13F,8'h06};
                12'd236  :cmd_data={1'b1,10'h13C,8'h00};
                12'd237  :cmd_data={1'b1,10'h13C,8'h00};
                12'd238  :cmd_data={1'b1,10'h13F,8'h02};
                12'd239  :cmd_data={1'b1,10'h13C,8'h00};
                12'd240  :cmd_data={1'b1,10'h13C,8'h00};
                12'd241  :cmd_data={1'b1,10'h13F,8'h00};
                12'd242  :cmd_data={1'b1,10'h137,8'h1A};
                12'd243  :cmd_data={1'b1,10'h130,8'h00};
                12'd244  :cmd_data={1'b1,10'h131,8'h00};
                12'd245  :cmd_data={1'b1,10'h132,8'h00};
                12'd246  :cmd_data={1'b1,10'h133,8'h20};
                12'd247  :cmd_data={1'b1,10'h137,8'h1E};
                12'd248  :cmd_data={1'b1,10'h134,8'h00};
                12'd249  :cmd_data={1'b1,10'h134,8'h00};
                12'd250  :cmd_data={1'b1,10'h130,8'h01};
                12'd251  :cmd_data={1'b1,10'h131,8'h00};
                12'd252  :cmd_data={1'b1,10'h132,8'h00};
                12'd253  :cmd_data={1'b1,10'h133,8'h00};
                12'd254  :cmd_data={1'b1,10'h137,8'h1E};
                12'd255  :cmd_data={1'b1,10'h134,8'h00};
                12'd256  :cmd_data={1'b1,10'h134,8'h00};
                12'd257  :cmd_data={1'b1,10'h130,8'h02};
                12'd258  :cmd_data={1'b1,10'h131,8'h00};
                12'd259  :cmd_data={1'b1,10'h132,8'h00};
                12'd260  :cmd_data={1'b1,10'h133,8'h00};
                12'd261  :cmd_data={1'b1,10'h137,8'h1E};
                12'd262  :cmd_data={1'b1,10'h134,8'h00};
                12'd263  :cmd_data={1'b1,10'h134,8'h00};
                12'd264  :cmd_data={1'b1,10'h130,8'h03};
                12'd265  :cmd_data={1'b1,10'h131,8'h00};
                12'd266  :cmd_data={1'b1,10'h132,8'h01};
                12'd267  :cmd_data={1'b1,10'h133,8'h00};
                12'd268  :cmd_data={1'b1,10'h137,8'h1E};
                12'd269  :cmd_data={1'b1,10'h134,8'h00};
                12'd270  :cmd_data={1'b1,10'h134,8'h00};
                12'd271  :cmd_data={1'b1,10'h130,8'h04};
                12'd272  :cmd_data={1'b1,10'h131,8'h00};
                12'd273  :cmd_data={1'b1,10'h132,8'h02};
                12'd274  :cmd_data={1'b1,10'h133,8'h00};
                12'd275  :cmd_data={1'b1,10'h137,8'h1E};
                12'd276  :cmd_data={1'b1,10'h134,8'h00};
                12'd277  :cmd_data={1'b1,10'h134,8'h00};
                12'd278  :cmd_data={1'b1,10'h130,8'h05};
                12'd279  :cmd_data={1'b1,10'h131,8'h00};
                12'd280  :cmd_data={1'b1,10'h132,8'h03};
                12'd281  :cmd_data={1'b1,10'h133,8'h00};
                12'd282  :cmd_data={1'b1,10'h137,8'h1E};
                12'd283  :cmd_data={1'b1,10'h134,8'h00};
                12'd284  :cmd_data={1'b1,10'h134,8'h00};
                12'd285  :cmd_data={1'b1,10'h130,8'h06};
                12'd286  :cmd_data={1'b1,10'h131,8'h00};
                12'd287  :cmd_data={1'b1,10'h132,8'h04};
                12'd288  :cmd_data={1'b1,10'h133,8'h00};
                12'd289  :cmd_data={1'b1,10'h137,8'h1E};
                12'd290  :cmd_data={1'b1,10'h134,8'h00};
                12'd291  :cmd_data={1'b1,10'h134,8'h00};
                12'd292  :cmd_data={1'b1,10'h130,8'h07};
                12'd293  :cmd_data={1'b1,10'h131,8'h00};
                12'd294  :cmd_data={1'b1,10'h132,8'h05};
                12'd295  :cmd_data={1'b1,10'h133,8'h00};
                12'd296  :cmd_data={1'b1,10'h137,8'h1E};
                12'd297  :cmd_data={1'b1,10'h134,8'h00};
                12'd298  :cmd_data={1'b1,10'h134,8'h00};
                12'd299  :cmd_data={1'b1,10'h130,8'h08};
                12'd300  :cmd_data={1'b1,10'h131,8'h01};
                12'd301  :cmd_data={1'b1,10'h132,8'h03};
                12'd302  :cmd_data={1'b1,10'h133,8'h20};
                12'd303  :cmd_data={1'b1,10'h137,8'h1E};
                12'd304  :cmd_data={1'b1,10'h134,8'h00};
                12'd305  :cmd_data={1'b1,10'h134,8'h00};
                12'd306  :cmd_data={1'b1,10'h130,8'h09};
                12'd307  :cmd_data={1'b1,10'h131,8'h01};
                12'd308  :cmd_data={1'b1,10'h132,8'h04};
                12'd309  :cmd_data={1'b1,10'h133,8'h00};
                12'd310  :cmd_data={1'b1,10'h137,8'h1E};
                12'd311  :cmd_data={1'b1,10'h134,8'h00};
                12'd312  :cmd_data={1'b1,10'h134,8'h00};
                12'd313  :cmd_data={1'b1,10'h130,8'h0A};
                12'd314  :cmd_data={1'b1,10'h131,8'h01};
                12'd315  :cmd_data={1'b1,10'h132,8'h05};
                12'd316  :cmd_data={1'b1,10'h133,8'h00};
                12'd317  :cmd_data={1'b1,10'h137,8'h1E};
                12'd318  :cmd_data={1'b1,10'h134,8'h00};
                12'd319  :cmd_data={1'b1,10'h134,8'h00};
                12'd320  :cmd_data={1'b1,10'h130,8'h0B};
                12'd321  :cmd_data={1'b1,10'h131,8'h01};
                12'd322  :cmd_data={1'b1,10'h132,8'h06};
                12'd323  :cmd_data={1'b1,10'h133,8'h00};
                12'd324  :cmd_data={1'b1,10'h137,8'h1E};
                12'd325  :cmd_data={1'b1,10'h134,8'h00};
                12'd326  :cmd_data={1'b1,10'h134,8'h00};
                12'd327  :cmd_data={1'b1,10'h130,8'h0C};
                12'd328  :cmd_data={1'b1,10'h131,8'h01};
                12'd329  :cmd_data={1'b1,10'h132,8'h07};
                12'd330  :cmd_data={1'b1,10'h133,8'h00};
                12'd331  :cmd_data={1'b1,10'h137,8'h1E};
                12'd332  :cmd_data={1'b1,10'h134,8'h00};
                12'd333  :cmd_data={1'b1,10'h134,8'h00};
                12'd334  :cmd_data={1'b1,10'h130,8'h0D};
                12'd335  :cmd_data={1'b1,10'h131,8'h01};
                12'd336  :cmd_data={1'b1,10'h132,8'h08};
                12'd337  :cmd_data={1'b1,10'h133,8'h00};
                12'd338  :cmd_data={1'b1,10'h137,8'h1E};
                12'd339  :cmd_data={1'b1,10'h134,8'h00};
                12'd340  :cmd_data={1'b1,10'h134,8'h00};
                12'd341  :cmd_data={1'b1,10'h130,8'h0E};
                12'd342  :cmd_data={1'b1,10'h131,8'h01};
                12'd343  :cmd_data={1'b1,10'h132,8'h09};
                12'd344  :cmd_data={1'b1,10'h133,8'h00};
                12'd345  :cmd_data={1'b1,10'h137,8'h1E};
                12'd346  :cmd_data={1'b1,10'h134,8'h00};
                12'd347  :cmd_data={1'b1,10'h134,8'h00};
                12'd348  :cmd_data={1'b1,10'h130,8'h0F};
                12'd349  :cmd_data={1'b1,10'h131,8'h01};
                12'd350  :cmd_data={1'b1,10'h132,8'h0A};
                12'd351  :cmd_data={1'b1,10'h133,8'h00};
                12'd352  :cmd_data={1'b1,10'h137,8'h1E};
                12'd353  :cmd_data={1'b1,10'h134,8'h00};
                12'd354  :cmd_data={1'b1,10'h134,8'h00};
                12'd355  :cmd_data={1'b1,10'h130,8'h10};
                12'd356  :cmd_data={1'b1,10'h131,8'h01};
                12'd357  :cmd_data={1'b1,10'h132,8'h0B};
                12'd358  :cmd_data={1'b1,10'h133,8'h00};
                12'd359  :cmd_data={1'b1,10'h137,8'h1E};
                12'd360  :cmd_data={1'b1,10'h134,8'h00};
                12'd361  :cmd_data={1'b1,10'h134,8'h00};
                12'd362  :cmd_data={1'b1,10'h130,8'h11};
                12'd363  :cmd_data={1'b1,10'h131,8'h01};
                12'd364  :cmd_data={1'b1,10'h132,8'h0C};
                12'd365  :cmd_data={1'b1,10'h133,8'h00};
                12'd366  :cmd_data={1'b1,10'h137,8'h1E};
                12'd367  :cmd_data={1'b1,10'h134,8'h00};
                12'd368  :cmd_data={1'b1,10'h134,8'h00};
                12'd369  :cmd_data={1'b1,10'h130,8'h12};
                12'd370  :cmd_data={1'b1,10'h131,8'h01};
                12'd371  :cmd_data={1'b1,10'h132,8'h0D};
                12'd372  :cmd_data={1'b1,10'h133,8'h00};
                12'd373  :cmd_data={1'b1,10'h137,8'h1E};
                12'd374  :cmd_data={1'b1,10'h134,8'h00};
                12'd375  :cmd_data={1'b1,10'h134,8'h00};
                12'd376  :cmd_data={1'b1,10'h130,8'h13};
                12'd377  :cmd_data={1'b1,10'h131,8'h01};
                12'd378  :cmd_data={1'b1,10'h132,8'h0E};
                12'd379  :cmd_data={1'b1,10'h133,8'h00};
                12'd380  :cmd_data={1'b1,10'h137,8'h1E};
                12'd381  :cmd_data={1'b1,10'h134,8'h00};
                12'd382  :cmd_data={1'b1,10'h134,8'h00};
                12'd383  :cmd_data={1'b1,10'h130,8'h14};
                12'd384  :cmd_data={1'b1,10'h131,8'h02};
                12'd385  :cmd_data={1'b1,10'h132,8'h09};
                12'd386  :cmd_data={1'b1,10'h133,8'h20};
                12'd387  :cmd_data={1'b1,10'h137,8'h1E};
                12'd388  :cmd_data={1'b1,10'h134,8'h00};
                12'd389  :cmd_data={1'b1,10'h134,8'h00};
                12'd390  :cmd_data={1'b1,10'h130,8'h15};
                12'd391  :cmd_data={1'b1,10'h131,8'h02};
                12'd392  :cmd_data={1'b1,10'h132,8'h0A};
                12'd393  :cmd_data={1'b1,10'h133,8'h00};
                12'd394  :cmd_data={1'b1,10'h137,8'h1E};
                12'd395  :cmd_data={1'b1,10'h134,8'h00};
                12'd396  :cmd_data={1'b1,10'h134,8'h00};
                12'd397  :cmd_data={1'b1,10'h130,8'h16};
                12'd398  :cmd_data={1'b1,10'h131,8'h02};
                12'd399  :cmd_data={1'b1,10'h132,8'h0B};
                12'd400  :cmd_data={1'b1,10'h133,8'h00};
                12'd401  :cmd_data={1'b1,10'h137,8'h1E};
                12'd402  :cmd_data={1'b1,10'h134,8'h00};
                12'd403  :cmd_data={1'b1,10'h134,8'h00};
                12'd404  :cmd_data={1'b1,10'h130,8'h17};
                12'd405  :cmd_data={1'b1,10'h131,8'h02};
                12'd406  :cmd_data={1'b1,10'h132,8'h0C};
                12'd407  :cmd_data={1'b1,10'h133,8'h00};
                12'd408  :cmd_data={1'b1,10'h137,8'h1E};
                12'd409  :cmd_data={1'b1,10'h134,8'h00};
                12'd410  :cmd_data={1'b1,10'h134,8'h00};
                12'd411  :cmd_data={1'b1,10'h130,8'h18};
                12'd412  :cmd_data={1'b1,10'h131,8'h02};
                12'd413  :cmd_data={1'b1,10'h132,8'h0D};
                12'd414  :cmd_data={1'b1,10'h133,8'h00};
                12'd415  :cmd_data={1'b1,10'h137,8'h1E};
                12'd416  :cmd_data={1'b1,10'h134,8'h00};
                12'd417  :cmd_data={1'b1,10'h134,8'h00};
                12'd418  :cmd_data={1'b1,10'h130,8'h19};
                12'd419  :cmd_data={1'b1,10'h131,8'h02};
                12'd420  :cmd_data={1'b1,10'h132,8'h0E};
                12'd421  :cmd_data={1'b1,10'h133,8'h00};
                12'd422  :cmd_data={1'b1,10'h137,8'h1E};
                12'd423  :cmd_data={1'b1,10'h134,8'h00};
                12'd424  :cmd_data={1'b1,10'h134,8'h00};
                12'd425  :cmd_data={1'b1,10'h130,8'h1A};
                12'd426  :cmd_data={1'b1,10'h131,8'h02};
                12'd427  :cmd_data={1'b1,10'h132,8'h0F};
                12'd428  :cmd_data={1'b1,10'h133,8'h00};
                12'd429  :cmd_data={1'b1,10'h137,8'h1E};
                12'd430  :cmd_data={1'b1,10'h134,8'h00};
                12'd431  :cmd_data={1'b1,10'h134,8'h00};
                12'd432  :cmd_data={1'b1,10'h130,8'h1B};
                12'd433  :cmd_data={1'b1,10'h131,8'h02};
                12'd434  :cmd_data={1'b1,10'h132,8'h10};
                12'd435  :cmd_data={1'b1,10'h133,8'h00};
                12'd436  :cmd_data={1'b1,10'h137,8'h1E};
                12'd437  :cmd_data={1'b1,10'h134,8'h00};
                12'd438  :cmd_data={1'b1,10'h134,8'h00};
                12'd439  :cmd_data={1'b1,10'h130,8'h1C};
                12'd440  :cmd_data={1'b1,10'h131,8'h02};
                12'd441  :cmd_data={1'b1,10'h132,8'h2B};
                12'd442  :cmd_data={1'b1,10'h133,8'h20};
                12'd443  :cmd_data={1'b1,10'h137,8'h1E};
                12'd444  :cmd_data={1'b1,10'h134,8'h00};
                12'd445  :cmd_data={1'b1,10'h134,8'h00};
                12'd446  :cmd_data={1'b1,10'h130,8'h1D};
                12'd447  :cmd_data={1'b1,10'h131,8'h02};
                12'd448  :cmd_data={1'b1,10'h132,8'h2C};
                12'd449  :cmd_data={1'b1,10'h133,8'h00};
                12'd450  :cmd_data={1'b1,10'h137,8'h1E};
                12'd451  :cmd_data={1'b1,10'h134,8'h00};
                12'd452  :cmd_data={1'b1,10'h134,8'h00};
                12'd453  :cmd_data={1'b1,10'h130,8'h1E};
                12'd454  :cmd_data={1'b1,10'h131,8'h04};
                12'd455  :cmd_data={1'b1,10'h132,8'h27};
                12'd456  :cmd_data={1'b1,10'h133,8'h20};
                12'd457  :cmd_data={1'b1,10'h137,8'h1E};
                12'd458  :cmd_data={1'b1,10'h134,8'h00};
                12'd459  :cmd_data={1'b1,10'h134,8'h00};
                12'd460  :cmd_data={1'b1,10'h130,8'h1F};
                12'd461  :cmd_data={1'b1,10'h131,8'h04};
                12'd462  :cmd_data={1'b1,10'h132,8'h28};
                12'd463  :cmd_data={1'b1,10'h133,8'h00};
                12'd464  :cmd_data={1'b1,10'h137,8'h1E};
                12'd465  :cmd_data={1'b1,10'h134,8'h00};
                12'd466  :cmd_data={1'b1,10'h134,8'h00};
                12'd467  :cmd_data={1'b1,10'h130,8'h20};
                12'd468  :cmd_data={1'b1,10'h131,8'h04};
                12'd469  :cmd_data={1'b1,10'h132,8'h29};
                12'd470  :cmd_data={1'b1,10'h133,8'h00};
                12'd471  :cmd_data={1'b1,10'h137,8'h1E};
                12'd472  :cmd_data={1'b1,10'h134,8'h00};
                12'd473  :cmd_data={1'b1,10'h134,8'h00};
                12'd474  :cmd_data={1'b1,10'h130,8'h21};
                12'd475  :cmd_data={1'b1,10'h131,8'h04};
                12'd476  :cmd_data={1'b1,10'h132,8'h2A};
                12'd477  :cmd_data={1'b1,10'h133,8'h00};
                12'd478  :cmd_data={1'b1,10'h137,8'h1E};
                12'd479  :cmd_data={1'b1,10'h134,8'h00};
                12'd480  :cmd_data={1'b1,10'h134,8'h00};
                12'd481  :cmd_data={1'b1,10'h130,8'h22};
                12'd482  :cmd_data={1'b1,10'h131,8'h04};
                12'd483  :cmd_data={1'b1,10'h132,8'h2B};
                12'd484  :cmd_data={1'b1,10'h133,8'h00};
                12'd485  :cmd_data={1'b1,10'h137,8'h1E};
                12'd486  :cmd_data={1'b1,10'h134,8'h00};
                12'd487  :cmd_data={1'b1,10'h134,8'h00};
                12'd488  :cmd_data={1'b1,10'h130,8'h23};
                12'd489  :cmd_data={1'b1,10'h131,8'h24};
                12'd490  :cmd_data={1'b1,10'h132,8'h21};
                12'd491  :cmd_data={1'b1,10'h133,8'h20};
                12'd492  :cmd_data={1'b1,10'h137,8'h1E};
                12'd493  :cmd_data={1'b1,10'h134,8'h00};
                12'd494  :cmd_data={1'b1,10'h134,8'h00};
                12'd495  :cmd_data={1'b1,10'h130,8'h24};
                12'd496  :cmd_data={1'b1,10'h131,8'h24};
                12'd497  :cmd_data={1'b1,10'h132,8'h22};
                12'd498  :cmd_data={1'b1,10'h133,8'h00};
                12'd499  :cmd_data={1'b1,10'h137,8'h1E};
                12'd500  :cmd_data={1'b1,10'h134,8'h00};
                12'd501  :cmd_data={1'b1,10'h134,8'h00};
                12'd502  :cmd_data={1'b1,10'h130,8'h25};
                12'd503  :cmd_data={1'b1,10'h131,8'h44};
                12'd504  :cmd_data={1'b1,10'h132,8'h20};
                12'd505  :cmd_data={1'b1,10'h133,8'h20};
                12'd506  :cmd_data={1'b1,10'h137,8'h1E};
                12'd507  :cmd_data={1'b1,10'h134,8'h00};
                12'd508  :cmd_data={1'b1,10'h134,8'h00};
                12'd509  :cmd_data={1'b1,10'h130,8'h26};
                12'd510  :cmd_data={1'b1,10'h131,8'h44};
                12'd511  :cmd_data={1'b1,10'h132,8'h21};
                12'd512  :cmd_data={1'b1,10'h133,8'h00};
                12'd513  :cmd_data={1'b1,10'h137,8'h1E};
                12'd514  :cmd_data={1'b1,10'h134,8'h00};
                12'd515  :cmd_data={1'b1,10'h134,8'h00};
                12'd516  :cmd_data={1'b1,10'h130,8'h27};
                12'd517  :cmd_data={1'b1,10'h131,8'h44};
                12'd518  :cmd_data={1'b1,10'h132,8'h22};
                12'd519  :cmd_data={1'b1,10'h133,8'h00};
                12'd520  :cmd_data={1'b1,10'h137,8'h1E};
                12'd521  :cmd_data={1'b1,10'h134,8'h00};
                12'd522  :cmd_data={1'b1,10'h134,8'h00};
                12'd523  :cmd_data={1'b1,10'h130,8'h28};
                12'd524  :cmd_data={1'b1,10'h131,8'h44};
                12'd525  :cmd_data={1'b1,10'h132,8'h23};
                12'd526  :cmd_data={1'b1,10'h133,8'h00};
                12'd527  :cmd_data={1'b1,10'h137,8'h1E};
                12'd528  :cmd_data={1'b1,10'h134,8'h00};
                12'd529  :cmd_data={1'b1,10'h134,8'h00};
                12'd530  :cmd_data={1'b1,10'h130,8'h29};
                12'd531  :cmd_data={1'b1,10'h131,8'h44};
                12'd532  :cmd_data={1'b1,10'h132,8'h24};
                12'd533  :cmd_data={1'b1,10'h133,8'h00};
                12'd534  :cmd_data={1'b1,10'h137,8'h1E};
                12'd535  :cmd_data={1'b1,10'h134,8'h00};
                12'd536  :cmd_data={1'b1,10'h134,8'h00};
                12'd537  :cmd_data={1'b1,10'h130,8'h2A};
                12'd538  :cmd_data={1'b1,10'h131,8'h44};
                12'd539  :cmd_data={1'b1,10'h132,8'h25};
                12'd540  :cmd_data={1'b1,10'h133,8'h00};
                12'd541  :cmd_data={1'b1,10'h137,8'h1E};
                12'd542  :cmd_data={1'b1,10'h134,8'h00};
                12'd543  :cmd_data={1'b1,10'h134,8'h00};
                12'd544  :cmd_data={1'b1,10'h130,8'h2B};
                12'd545  :cmd_data={1'b1,10'h131,8'h44};
                12'd546  :cmd_data={1'b1,10'h132,8'h26};
                12'd547  :cmd_data={1'b1,10'h133,8'h00};
                12'd548  :cmd_data={1'b1,10'h137,8'h1E};
                12'd549  :cmd_data={1'b1,10'h134,8'h00};
                12'd550  :cmd_data={1'b1,10'h134,8'h00};
                12'd551  :cmd_data={1'b1,10'h130,8'h2C};
                12'd552  :cmd_data={1'b1,10'h131,8'h44};
                12'd553  :cmd_data={1'b1,10'h132,8'h27};
                12'd554  :cmd_data={1'b1,10'h133,8'h00};
                12'd555  :cmd_data={1'b1,10'h137,8'h1E};
                12'd556  :cmd_data={1'b1,10'h134,8'h00};
                12'd557  :cmd_data={1'b1,10'h134,8'h00};
                12'd558  :cmd_data={1'b1,10'h130,8'h2D};
                12'd559  :cmd_data={1'b1,10'h131,8'h44};
                12'd560  :cmd_data={1'b1,10'h132,8'h28};
                12'd561  :cmd_data={1'b1,10'h133,8'h00};
                12'd562  :cmd_data={1'b1,10'h137,8'h1E};
                12'd563  :cmd_data={1'b1,10'h134,8'h00};
                12'd564  :cmd_data={1'b1,10'h134,8'h00};
                12'd565  :cmd_data={1'b1,10'h130,8'h2E};
                12'd566  :cmd_data={1'b1,10'h131,8'h44};
                12'd567  :cmd_data={1'b1,10'h132,8'h29};
                12'd568  :cmd_data={1'b1,10'h133,8'h00};
                12'd569  :cmd_data={1'b1,10'h137,8'h1E};
                12'd570  :cmd_data={1'b1,10'h134,8'h00};
                12'd571  :cmd_data={1'b1,10'h134,8'h00};
                12'd572  :cmd_data={1'b1,10'h130,8'h2F};
                12'd573  :cmd_data={1'b1,10'h131,8'h44};
                12'd574  :cmd_data={1'b1,10'h132,8'h2A};
                12'd575  :cmd_data={1'b1,10'h133,8'h00};
                12'd576  :cmd_data={1'b1,10'h137,8'h1E};
                12'd577  :cmd_data={1'b1,10'h134,8'h00};
                12'd578  :cmd_data={1'b1,10'h134,8'h00};
                12'd579  :cmd_data={1'b1,10'h130,8'h30};
                12'd580  :cmd_data={1'b1,10'h131,8'h44};
                12'd581  :cmd_data={1'b1,10'h132,8'h2B};
                12'd582  :cmd_data={1'b1,10'h133,8'h00};
                12'd583  :cmd_data={1'b1,10'h137,8'h1E};
                12'd584  :cmd_data={1'b1,10'h134,8'h00};
                12'd585  :cmd_data={1'b1,10'h134,8'h00};
                12'd586  :cmd_data={1'b1,10'h130,8'h31};
                12'd587  :cmd_data={1'b1,10'h131,8'h44};
                12'd588  :cmd_data={1'b1,10'h132,8'h2C};
                12'd589  :cmd_data={1'b1,10'h133,8'h00};
                12'd590  :cmd_data={1'b1,10'h137,8'h1E};
                12'd591  :cmd_data={1'b1,10'h134,8'h00};
                12'd592  :cmd_data={1'b1,10'h134,8'h00};
                12'd593  :cmd_data={1'b1,10'h130,8'h32};
                12'd594  :cmd_data={1'b1,10'h131,8'h44};
                12'd595  :cmd_data={1'b1,10'h132,8'h2D};
                12'd596  :cmd_data={1'b1,10'h133,8'h00};
                12'd597  :cmd_data={1'b1,10'h137,8'h1E};
                12'd598  :cmd_data={1'b1,10'h134,8'h00};
                12'd599  :cmd_data={1'b1,10'h134,8'h00};
                12'd600  :cmd_data={1'b1,10'h130,8'h33};
                12'd601  :cmd_data={1'b1,10'h131,8'h44};
                12'd602  :cmd_data={1'b1,10'h132,8'h2E};
                12'd603  :cmd_data={1'b1,10'h133,8'h00};
                12'd604  :cmd_data={1'b1,10'h137,8'h1E};
                12'd605  :cmd_data={1'b1,10'h134,8'h00};
                12'd606  :cmd_data={1'b1,10'h134,8'h00};
                12'd607  :cmd_data={1'b1,10'h130,8'h34};
                12'd608  :cmd_data={1'b1,10'h131,8'h44};
                12'd609  :cmd_data={1'b1,10'h132,8'h2F};
                12'd610  :cmd_data={1'b1,10'h133,8'h00};
                12'd611  :cmd_data={1'b1,10'h137,8'h1E};
                12'd612  :cmd_data={1'b1,10'h134,8'h00};
                12'd613  :cmd_data={1'b1,10'h134,8'h00};
                12'd614  :cmd_data={1'b1,10'h130,8'h35};
                12'd615  :cmd_data={1'b1,10'h131,8'h44};
                12'd616  :cmd_data={1'b1,10'h132,8'h30};
                12'd617  :cmd_data={1'b1,10'h133,8'h00};
                12'd618  :cmd_data={1'b1,10'h137,8'h1E};
                12'd619  :cmd_data={1'b1,10'h134,8'h00};
                12'd620  :cmd_data={1'b1,10'h134,8'h00};
                12'd621  :cmd_data={1'b1,10'h130,8'h36};
                12'd622  :cmd_data={1'b1,10'h131,8'h44};
                12'd623  :cmd_data={1'b1,10'h132,8'h31};
                12'd624  :cmd_data={1'b1,10'h133,8'h00};
                12'd625  :cmd_data={1'b1,10'h137,8'h1E};
                12'd626  :cmd_data={1'b1,10'h134,8'h00};
                12'd627  :cmd_data={1'b1,10'h134,8'h00};
                12'd628  :cmd_data={1'b1,10'h130,8'h37};
                12'd629  :cmd_data={1'b1,10'h131,8'h64};
                12'd630  :cmd_data={1'b1,10'h132,8'h2E};
                12'd631  :cmd_data={1'b1,10'h133,8'h20};
                12'd632  :cmd_data={1'b1,10'h137,8'h1E};
                12'd633  :cmd_data={1'b1,10'h134,8'h00};
                12'd634  :cmd_data={1'b1,10'h134,8'h00};
                12'd635  :cmd_data={1'b1,10'h130,8'h38};
                12'd636  :cmd_data={1'b1,10'h131,8'h64};
                12'd637  :cmd_data={1'b1,10'h132,8'h2F};
                12'd638  :cmd_data={1'b1,10'h133,8'h00};
                12'd639  :cmd_data={1'b1,10'h137,8'h1E};
                12'd640  :cmd_data={1'b1,10'h134,8'h00};
                12'd641  :cmd_data={1'b1,10'h134,8'h00};
                12'd642  :cmd_data={1'b1,10'h130,8'h39};
                12'd643  :cmd_data={1'b1,10'h131,8'h64};
                12'd644  :cmd_data={1'b1,10'h132,8'h30};
                12'd645  :cmd_data={1'b1,10'h133,8'h00};
                12'd646  :cmd_data={1'b1,10'h137,8'h1E};
                12'd647  :cmd_data={1'b1,10'h134,8'h00};
                12'd648  :cmd_data={1'b1,10'h134,8'h00};
                12'd649  :cmd_data={1'b1,10'h130,8'h3A};
                12'd650  :cmd_data={1'b1,10'h131,8'h64};
                12'd651  :cmd_data={1'b1,10'h132,8'h31};
                12'd652  :cmd_data={1'b1,10'h133,8'h00};
                12'd653  :cmd_data={1'b1,10'h137,8'h1E};
                12'd654  :cmd_data={1'b1,10'h134,8'h00};
                12'd655  :cmd_data={1'b1,10'h134,8'h00};
                12'd656  :cmd_data={1'b1,10'h130,8'h3B};
                12'd657  :cmd_data={1'b1,10'h131,8'h64};
                12'd658  :cmd_data={1'b1,10'h132,8'h32};
                12'd659  :cmd_data={1'b1,10'h133,8'h00};
                12'd660  :cmd_data={1'b1,10'h137,8'h1E};
                12'd661  :cmd_data={1'b1,10'h134,8'h00};
                12'd662  :cmd_data={1'b1,10'h134,8'h00};
                12'd663  :cmd_data={1'b1,10'h130,8'h3C};
                12'd664  :cmd_data={1'b1,10'h131,8'h64};
                12'd665  :cmd_data={1'b1,10'h132,8'h33};
                12'd666  :cmd_data={1'b1,10'h133,8'h00};
                12'd667  :cmd_data={1'b1,10'h137,8'h1E};
                12'd668  :cmd_data={1'b1,10'h134,8'h00};
                12'd669  :cmd_data={1'b1,10'h134,8'h00};
                12'd670  :cmd_data={1'b1,10'h130,8'h3D};
                12'd671  :cmd_data={1'b1,10'h131,8'h64};
                12'd672  :cmd_data={1'b1,10'h132,8'h34};
                12'd673  :cmd_data={1'b1,10'h133,8'h00};
                12'd674  :cmd_data={1'b1,10'h137,8'h1E};
                12'd675  :cmd_data={1'b1,10'h134,8'h00};
                12'd676  :cmd_data={1'b1,10'h134,8'h00};
                12'd677  :cmd_data={1'b1,10'h130,8'h3E};
                12'd678  :cmd_data={1'b1,10'h131,8'h64};
                12'd679  :cmd_data={1'b1,10'h132,8'h35};
                12'd680  :cmd_data={1'b1,10'h133,8'h00};
                12'd681  :cmd_data={1'b1,10'h137,8'h1E};
                12'd682  :cmd_data={1'b1,10'h134,8'h00};
                12'd683  :cmd_data={1'b1,10'h134,8'h00};
                12'd684  :cmd_data={1'b1,10'h130,8'h3F};
                12'd685  :cmd_data={1'b1,10'h131,8'h64};
                12'd686  :cmd_data={1'b1,10'h132,8'h36};
                12'd687  :cmd_data={1'b1,10'h133,8'h00};
                12'd688  :cmd_data={1'b1,10'h137,8'h1E};
                12'd689  :cmd_data={1'b1,10'h134,8'h00};
                12'd690  :cmd_data={1'b1,10'h134,8'h00};
                12'd691  :cmd_data={1'b1,10'h130,8'h40};
                12'd692  :cmd_data={1'b1,10'h131,8'h64};
                12'd693  :cmd_data={1'b1,10'h132,8'h37};
                12'd694  :cmd_data={1'b1,10'h133,8'h00};
                12'd695  :cmd_data={1'b1,10'h137,8'h1E};
                12'd696  :cmd_data={1'b1,10'h134,8'h00};
                12'd697  :cmd_data={1'b1,10'h134,8'h00};
                12'd698  :cmd_data={1'b1,10'h130,8'h41};
                12'd699  :cmd_data={1'b1,10'h131,8'h64};
                12'd700  :cmd_data={1'b1,10'h132,8'h38};
                12'd701  :cmd_data={1'b1,10'h133,8'h00};
                12'd702  :cmd_data={1'b1,10'h137,8'h1E};
                12'd703  :cmd_data={1'b1,10'h134,8'h00};
                12'd704  :cmd_data={1'b1,10'h134,8'h00};
                12'd705  :cmd_data={1'b1,10'h130,8'h42};
                12'd706  :cmd_data={1'b1,10'h131,8'h65};
                12'd707  :cmd_data={1'b1,10'h132,8'h38};
                12'd708  :cmd_data={1'b1,10'h133,8'h20};
                12'd709  :cmd_data={1'b1,10'h137,8'h1E};
                12'd710  :cmd_data={1'b1,10'h134,8'h00};
                12'd711  :cmd_data={1'b1,10'h134,8'h00};
                12'd712  :cmd_data={1'b1,10'h130,8'h43};
                12'd713  :cmd_data={1'b1,10'h131,8'h66};
                12'd714  :cmd_data={1'b1,10'h132,8'h38};
                12'd715  :cmd_data={1'b1,10'h133,8'h20};
                12'd716  :cmd_data={1'b1,10'h137,8'h1E};
                12'd717  :cmd_data={1'b1,10'h134,8'h00};
                12'd718  :cmd_data={1'b1,10'h134,8'h00};
                12'd719  :cmd_data={1'b1,10'h130,8'h44};
                12'd720  :cmd_data={1'b1,10'h131,8'h67};
                12'd721  :cmd_data={1'b1,10'h132,8'h38};
                12'd722  :cmd_data={1'b1,10'h133,8'h20};
                12'd723  :cmd_data={1'b1,10'h137,8'h1E};
                12'd724  :cmd_data={1'b1,10'h134,8'h00};
                12'd725  :cmd_data={1'b1,10'h134,8'h00};
                12'd726  :cmd_data={1'b1,10'h130,8'h45};
                12'd727  :cmd_data={1'b1,10'h131,8'h68};
                12'd728  :cmd_data={1'b1,10'h132,8'h38};
                12'd729  :cmd_data={1'b1,10'h133,8'h20};
                12'd730  :cmd_data={1'b1,10'h137,8'h1E};
                12'd731  :cmd_data={1'b1,10'h134,8'h00};
                12'd732  :cmd_data={1'b1,10'h134,8'h00};
                12'd733  :cmd_data={1'b1,10'h130,8'h46};
                12'd734  :cmd_data={1'b1,10'h131,8'h69};
                12'd735  :cmd_data={1'b1,10'h132,8'h38};
                12'd736  :cmd_data={1'b1,10'h133,8'h20};
                12'd737  :cmd_data={1'b1,10'h137,8'h1E};
                12'd738  :cmd_data={1'b1,10'h134,8'h00};
                12'd739  :cmd_data={1'b1,10'h134,8'h00};
                12'd740  :cmd_data={1'b1,10'h130,8'h47};
                12'd741  :cmd_data={1'b1,10'h131,8'h6A};
                12'd742  :cmd_data={1'b1,10'h132,8'h38};
                12'd743  :cmd_data={1'b1,10'h133,8'h20};
                12'd744  :cmd_data={1'b1,10'h137,8'h1E};
                12'd745  :cmd_data={1'b1,10'h134,8'h00};
                12'd746  :cmd_data={1'b1,10'h134,8'h00};
                12'd747  :cmd_data={1'b1,10'h130,8'h48};
                12'd748  :cmd_data={1'b1,10'h131,8'h6B};
                12'd749  :cmd_data={1'b1,10'h132,8'h38};
                12'd750  :cmd_data={1'b1,10'h133,8'h20};
                12'd751  :cmd_data={1'b1,10'h137,8'h1E};
                12'd752  :cmd_data={1'b1,10'h134,8'h00};
                12'd753  :cmd_data={1'b1,10'h134,8'h00};
                12'd754  :cmd_data={1'b1,10'h130,8'h49};
                12'd755  :cmd_data={1'b1,10'h131,8'h6C};
                12'd756  :cmd_data={1'b1,10'h132,8'h38};
                12'd757  :cmd_data={1'b1,10'h133,8'h20};
                12'd758  :cmd_data={1'b1,10'h137,8'h1E};
                12'd759  :cmd_data={1'b1,10'h134,8'h00};
                12'd760  :cmd_data={1'b1,10'h134,8'h00};
                12'd761  :cmd_data={1'b1,10'h130,8'h4A};
                12'd762  :cmd_data={1'b1,10'h131,8'h6D};
                12'd763  :cmd_data={1'b1,10'h132,8'h38};
                12'd764  :cmd_data={1'b1,10'h133,8'h20};
                12'd765  :cmd_data={1'b1,10'h137,8'h1E};
                12'd766  :cmd_data={1'b1,10'h134,8'h00};
                12'd767  :cmd_data={1'b1,10'h134,8'h00};
                12'd768  :cmd_data={1'b1,10'h130,8'h4B};
                12'd769  :cmd_data={1'b1,10'h131,8'h6E};
                12'd770  :cmd_data={1'b1,10'h132,8'h38};
                12'd771  :cmd_data={1'b1,10'h133,8'h20};
                12'd772  :cmd_data={1'b1,10'h137,8'h1E};
                12'd773  :cmd_data={1'b1,10'h134,8'h00};
                12'd774  :cmd_data={1'b1,10'h134,8'h00};
                12'd775  :cmd_data={1'b1,10'h130,8'h4C};
                12'd776  :cmd_data={1'b1,10'h131,8'h6F};
                12'd777  :cmd_data={1'b1,10'h132,8'h38};
                12'd778  :cmd_data={1'b1,10'h133,8'h20};
                12'd779  :cmd_data={1'b1,10'h137,8'h1E};
                12'd780  :cmd_data={1'b1,10'h134,8'h00};
                12'd781  :cmd_data={1'b1,10'h134,8'h00};
                12'd782  :cmd_data={1'b1,10'h130,8'h4D};
                12'd783  :cmd_data={1'b1,10'h131,8'h00};
                12'd784  :cmd_data={1'b1,10'h132,8'h00};
                12'd785  :cmd_data={1'b1,10'h133,8'h00};
                12'd786  :cmd_data={1'b1,10'h137,8'h1E};
                12'd787  :cmd_data={1'b1,10'h134,8'h00};
                12'd788  :cmd_data={1'b1,10'h134,8'h00};
                12'd789  :cmd_data={1'b1,10'h130,8'h4E};
                12'd790  :cmd_data={1'b1,10'h131,8'h00};
                12'd791  :cmd_data={1'b1,10'h132,8'h00};
                12'd792  :cmd_data={1'b1,10'h133,8'h00};
                12'd793  :cmd_data={1'b1,10'h137,8'h1E};
                12'd794  :cmd_data={1'b1,10'h134,8'h00};
                12'd795  :cmd_data={1'b1,10'h134,8'h00};
                12'd796  :cmd_data={1'b1,10'h130,8'h4F};
                12'd797  :cmd_data={1'b1,10'h131,8'h00};
                12'd798  :cmd_data={1'b1,10'h132,8'h00};
                12'd799  :cmd_data={1'b1,10'h133,8'h00};
                12'd800  :cmd_data={1'b1,10'h137,8'h1E};
                12'd801  :cmd_data={1'b1,10'h134,8'h00};
                12'd802  :cmd_data={1'b1,10'h134,8'h00};
                12'd803  :cmd_data={1'b1,10'h130,8'h50};
                12'd804  :cmd_data={1'b1,10'h131,8'h00};
                12'd805  :cmd_data={1'b1,10'h132,8'h00};
                12'd806  :cmd_data={1'b1,10'h133,8'h00};
                12'd807  :cmd_data={1'b1,10'h137,8'h1E};
                12'd808  :cmd_data={1'b1,10'h134,8'h00};
                12'd809  :cmd_data={1'b1,10'h134,8'h00};
                12'd810  :cmd_data={1'b1,10'h130,8'h51};
                12'd811  :cmd_data={1'b1,10'h131,8'h00};
                12'd812  :cmd_data={1'b1,10'h132,8'h00};
                12'd813  :cmd_data={1'b1,10'h133,8'h00};
                12'd814  :cmd_data={1'b1,10'h137,8'h1E};
                12'd815  :cmd_data={1'b1,10'h134,8'h00};
                12'd816  :cmd_data={1'b1,10'h134,8'h00};
                12'd817  :cmd_data={1'b1,10'h130,8'h52};
                12'd818  :cmd_data={1'b1,10'h131,8'h00};
                12'd819  :cmd_data={1'b1,10'h132,8'h00};
                12'd820  :cmd_data={1'b1,10'h133,8'h00};
                12'd821  :cmd_data={1'b1,10'h137,8'h1E};
                12'd822  :cmd_data={1'b1,10'h134,8'h00};
                12'd823  :cmd_data={1'b1,10'h134,8'h00};
                12'd824  :cmd_data={1'b1,10'h130,8'h53};
                12'd825  :cmd_data={1'b1,10'h131,8'h00};
                12'd826  :cmd_data={1'b1,10'h132,8'h00};
                12'd827  :cmd_data={1'b1,10'h133,8'h00};
                12'd828  :cmd_data={1'b1,10'h137,8'h1E};
                12'd829  :cmd_data={1'b1,10'h134,8'h00};
                12'd830  :cmd_data={1'b1,10'h134,8'h00};
                12'd831  :cmd_data={1'b1,10'h130,8'h54};
                12'd832  :cmd_data={1'b1,10'h131,8'h00};
                12'd833  :cmd_data={1'b1,10'h132,8'h00};
                12'd834  :cmd_data={1'b1,10'h133,8'h00};
                12'd835  :cmd_data={1'b1,10'h137,8'h1E};
                12'd836  :cmd_data={1'b1,10'h134,8'h00};
                12'd837  :cmd_data={1'b1,10'h134,8'h00};
                12'd838  :cmd_data={1'b1,10'h130,8'h55};
                12'd839  :cmd_data={1'b1,10'h131,8'h00};
                12'd840  :cmd_data={1'b1,10'h132,8'h00};
                12'd841  :cmd_data={1'b1,10'h133,8'h00};
                12'd842  :cmd_data={1'b1,10'h137,8'h1E};
                12'd843  :cmd_data={1'b1,10'h134,8'h00};
                12'd844  :cmd_data={1'b1,10'h134,8'h00};
                12'd845  :cmd_data={1'b1,10'h130,8'h56};
                12'd846  :cmd_data={1'b1,10'h131,8'h00};
                12'd847  :cmd_data={1'b1,10'h132,8'h00};
                12'd848  :cmd_data={1'b1,10'h133,8'h00};
                12'd849  :cmd_data={1'b1,10'h137,8'h1E};
                12'd850  :cmd_data={1'b1,10'h134,8'h00};
                12'd851  :cmd_data={1'b1,10'h134,8'h00};
                12'd852  :cmd_data={1'b1,10'h130,8'h57};
                12'd853  :cmd_data={1'b1,10'h131,8'h00};
                12'd854  :cmd_data={1'b1,10'h132,8'h00};
                12'd855  :cmd_data={1'b1,10'h133,8'h00};
                12'd856  :cmd_data={1'b1,10'h137,8'h1E};
                12'd857  :cmd_data={1'b1,10'h134,8'h00};
                12'd858  :cmd_data={1'b1,10'h134,8'h00};
                12'd859  :cmd_data={1'b1,10'h130,8'h58};
                12'd860  :cmd_data={1'b1,10'h131,8'h00};
                12'd861  :cmd_data={1'b1,10'h132,8'h00};
                12'd862  :cmd_data={1'b1,10'h133,8'h00};
                12'd863  :cmd_data={1'b1,10'h137,8'h1E};
                12'd864  :cmd_data={1'b1,10'h134,8'h00};
                12'd865  :cmd_data={1'b1,10'h134,8'h00};
                12'd866  :cmd_data={1'b1,10'h130,8'h59};
                12'd867  :cmd_data={1'b1,10'h131,8'h00};
                12'd868  :cmd_data={1'b1,10'h132,8'h00};
                12'd869  :cmd_data={1'b1,10'h133,8'h00};
                12'd870  :cmd_data={1'b1,10'h137,8'h1E};
                12'd871  :cmd_data={1'b1,10'h134,8'h00};
                12'd872  :cmd_data={1'b1,10'h134,8'h00};
                12'd873  :cmd_data={1'b1,10'h130,8'h5A};
                12'd874  :cmd_data={1'b1,10'h131,8'h00};
                12'd875  :cmd_data={1'b1,10'h132,8'h00};
                12'd876  :cmd_data={1'b1,10'h133,8'h00};
                12'd877  :cmd_data={1'b1,10'h137,8'h1E};
                12'd878  :cmd_data={1'b1,10'h134,8'h00};
                12'd879  :cmd_data={1'b1,10'h134,8'h00};
                12'd880  :cmd_data={1'b1,10'h137,8'h1A};
                12'd881  :cmd_data={1'b1,10'h134,8'h00};
                12'd882  :cmd_data={1'b1,10'h134,8'h00};
                12'd883  :cmd_data={1'b1,10'h137,8'h00};
                12'd884  :cmd_data={1'b1,10'h0FA,8'hE0};
                12'd885  :cmd_data={1'b1,10'h0FB,8'h08};
                12'd886  :cmd_data={1'b1,10'h0FC,8'h23};
                12'd887  :cmd_data={1'b1,10'h0FD,8'h4C};
                12'd888  :cmd_data={1'b1,10'h0FE,8'h44};
                12'd889  :cmd_data={1'b1,10'h100,8'h6F};
                12'd890  :cmd_data={1'b1,10'h104,8'h2F};
                12'd891  :cmd_data={1'b1,10'h105,8'h3A};
                12'd892  :cmd_data={1'b1,10'h107,8'h2B};
                12'd893  :cmd_data={1'b1,10'h108,8'h31};
                12'd894  :cmd_data={1'b1,10'h109,8'h4C};
                12'd895  :cmd_data={1'b1,10'h10A,8'h58};
                12'd896  :cmd_data={1'b1,10'h10B,8'h00};
                12'd897  :cmd_data={1'b1,10'h10C,8'h4C};
                12'd898  :cmd_data={1'b1,10'h10D,8'h18};
                12'd899  :cmd_data={1'b1,10'h10E,8'h00};
                12'd900  :cmd_data={1'b1,10'h114,8'h30};
                12'd901  :cmd_data={1'b1,10'h11A,8'h27};
                12'd902  :cmd_data={1'b1,10'h081,8'h00};
                12'd903  :cmd_data={1'b1,10'h1FB,8'h1C};
                12'd904  :cmd_data={1'b1,10'h1FC,8'h00};
                12'd905  :cmd_data={1'b1,10'h1F8,8'h03};
                12'd906  :cmd_data={1'b1,10'h1F9,8'h1E};
                12'd907  :cmd_data={1'b1,10'h1D5,8'h3F};
                12'd908  :cmd_data={1'b1,10'h1C0,8'h03};
                12'd909  :cmd_data={1'b1,10'h1E2,8'h02};
                12'd910  :cmd_data={1'b1,10'h1E3,8'h02};
                12'd911  :cmd_data={1'b1,10'h016,8'h80};
                12'd912  :cmd_data={1'b0,10'h016,8'h00};
                12'd913  :cmd_data={1'b1,10'h1E2,8'h03};
                12'd914  :cmd_data={1'b1,10'h1E3,8'h03};
                12'd915  :cmd_data={1'b1,10'h0D6,8'h03};
                12'd916  :cmd_data={1'b1,10'h0D7,8'h1E};
                12'd917  :cmd_data={1'b1,10'h0CA,8'h22};
                12'd918  :cmd_data={1'b1,10'h016,8'h40};
                12'd919  :cmd_data={1'b0,10'h016,8'h01};
                12'd920  :cmd_data={1'b1,10'h0CA,8'h26};
                12'd921  :cmd_data={1'b0,10'h1EB,8'h00};
                12'd922  :cmd_data={1'b0,10'h1EC,8'h00};
                12'd923  :cmd_data={1'b0,10'h1E6,8'h00};
                12'd924  :cmd_data={1'b1,10'h1DB,8'h20};
                12'd925  :cmd_data={1'b1,10'h1DD,8'h00};
                12'd926  :cmd_data={1'b1,10'h1DF,8'h00};
                12'd927  :cmd_data={1'b1,10'h1DC,8'h46};
                12'd928  :cmd_data={1'b1,10'h1DE,8'h46};
                12'd929  :cmd_data={1'b1,10'h0D2,8'h04};
                12'd930  :cmd_data={1'b1,10'h0D1,8'h0C};
                12'd931  :cmd_data={1'b1,10'h0D0,8'h57};
                12'd932  :cmd_data={1'b0,10'h1EB,8'h00};
                12'd933  :cmd_data={1'b0,10'h1EC,8'h00};
                12'd934  :cmd_data={1'b0,10'h1E6,8'h00};
                12'd935  :cmd_data={1'b1,10'h200,8'h00};
                12'd936  :cmd_data={1'b1,10'h201,8'h00};
                12'd937  :cmd_data={1'b1,10'h202,8'h00};
                12'd938  :cmd_data={1'b1,10'h203,8'h24};
                12'd939  :cmd_data={1'b1,10'h204,8'h24};
                12'd940  :cmd_data={1'b1,10'h205,8'h00};
                12'd941  :cmd_data={1'b1,10'h206,8'h00};
                12'd942  :cmd_data={1'b1,10'h207,8'h71};
                12'd943  :cmd_data={1'b1,10'h208,8'h71};
                12'd944  :cmd_data={1'b1,10'h209,8'h36};
                12'd945  :cmd_data={1'b1,10'h20A,8'h44};
                12'd946  :cmd_data={1'b1,10'h20B,8'h47};
                12'd947  :cmd_data={1'b1,10'h20C,8'h47};
                12'd948  :cmd_data={1'b1,10'h20D,8'h45};
                12'd949  :cmd_data={1'b1,10'h20E,8'h00};
                12'd950  :cmd_data={1'b1,10'h20F,8'h74};
                12'd951  :cmd_data={1'b1,10'h210,8'h74};
                12'd952  :cmd_data={1'b1,10'h211,8'h74};
                12'd953  :cmd_data={1'b1,10'h212,8'h42};
                12'd954  :cmd_data={1'b1,10'h213,8'h42};
                12'd955  :cmd_data={1'b1,10'h214,8'h42};
                12'd956  :cmd_data={1'b1,10'h215,8'h45};
                12'd957  :cmd_data={1'b1,10'h216,8'h45};
                12'd958  :cmd_data={1'b1,10'h217,8'h45};
                12'd959  :cmd_data={1'b1,10'h218,8'h2E};
                12'd960  :cmd_data={1'b1,10'h219,8'h93};
                12'd961  :cmd_data={1'b1,10'h21A,8'h17};
                12'd962  :cmd_data={1'b1,10'h21B,8'h11};
                12'd963  :cmd_data={1'b1,10'h21C,8'h93};
                12'd964  :cmd_data={1'b1,10'h21D,8'h17};
                12'd965  :cmd_data={1'b1,10'h21E,8'h11};
                12'd966  :cmd_data={1'b1,10'h21F,8'h93};
                12'd967  :cmd_data={1'b1,10'h220,8'h17};
                12'd968  :cmd_data={1'b1,10'h221,8'h23};
                12'd969  :cmd_data={1'b1,10'h222,8'h23};
                12'd970  :cmd_data={1'b1,10'h223,8'h40};
                12'd971  :cmd_data={1'b1,10'h224,8'h40};
                12'd972  :cmd_data={1'b1,10'h225,8'h2C};
                12'd973  :cmd_data={1'b1,10'h226,8'h00};
                12'd974  :cmd_data={1'b1,10'h227,8'h00};
                12'd975  :cmd_data={1'b1,10'h193,8'h3F};
                12'd976  :cmd_data={1'b1,10'h190,8'h0F};
                12'd977  :cmd_data={1'b1,10'h194,8'h01};
                12'd978  :cmd_data={1'b1,10'h016,8'h01};
                12'd979  :cmd_data={1'b0,10'h016,8'h02};
                12'd980  :cmd_data={1'b1,10'h185,8'h20};
                12'd981  :cmd_data={1'b1,10'h186,8'h32};
                12'd982  :cmd_data={1'b1,10'h187,8'h24};
                12'd983  :cmd_data={1'b1,10'h18B,8'h83};
                12'd984  :cmd_data={1'b1,10'h188,8'h05};
                12'd985  :cmd_data={1'b1,10'h189,8'h30};
                12'd986  :cmd_data={1'b1,10'h016,8'h02};
                12'd987  :cmd_data={1'b1,10'hFFF,8'hFF};
                12'd988  :cmd_data={1'b0,10'h0A3,8'h00};
                12'd989  :cmd_data={1'b1,10'h0A0,8'h3A};
                12'd990  :cmd_data={1'b1,10'h0A3,8'h40};
                12'd991  :cmd_data={1'b1,10'h0A1,8'h7B};
                12'd992  :cmd_data={1'b1,10'h0A9,8'hFF};
                12'd993  :cmd_data={1'b1,10'h0A2,8'h7F};
                12'd994  :cmd_data={1'b1,10'h0A5,8'h01};
                12'd995  :cmd_data={1'b1,10'h0A6,8'h01};
                12'd996  :cmd_data={1'b1,10'h0AA,8'h25};
                12'd997  :cmd_data={1'b1,10'h0A4,8'hF0};
                12'd998  :cmd_data={1'b1,10'h0AE,8'h00};
                12'd999  :cmd_data={1'b1,10'h169,8'hC0};
                12'd1000  :cmd_data={1'b1,10'h016,8'h10};
                12'd1001  :cmd_data={1'b0,10'h016,8'h03};
                12'd1002  :cmd_data={1'b1,10'h16A,8'h75};
                12'd1003  :cmd_data={1'b1,10'h16B,8'h95};
                12'd1004  :cmd_data={1'b1,10'h169,8'hCF};
                12'd1005  :cmd_data={1'b1,10'h18B,8'hAD};
                12'd1006  :cmd_data={1'b1,10'h012,8'h10};
                12'd1007  :cmd_data={1'b1,10'h013,8'h00};
                12'd1008  :cmd_data={1'b1,10'h015,8'h00};
                12'd1009  :cmd_data={1'b1,10'h073,8'h28};
                12'd1010  :cmd_data={1'b1,10'h074,8'h00};
                12'd1011  :cmd_data={1'b1,10'h075,8'h28};
                12'd1012  :cmd_data={1'b1,10'h076,8'h00};
                12'd1013  :cmd_data={1'b1,10'h150,8'h0E};
                12'd1014  :cmd_data={1'b1,10'h151,8'h00};
                12'd1015  :cmd_data={1'b1,10'h152,8'hFF};
                12'd1016  :cmd_data={1'b1,10'h153,8'h00};
                12'd1017  :cmd_data={1'b1,10'h154,8'h00};
                12'd1018  :cmd_data={1'b1,10'h155,8'h00};
                12'd1019  :cmd_data={1'b1,10'h156,8'h00};
                12'd1020  :cmd_data={1'b1,10'h157,8'h00};
                12'd1021  :cmd_data={1'b1,10'h158,8'h0D};
                12'd1022  :cmd_data={1'b1,10'h15C,8'h67};
                12'd1023  :cmd_data={1'b1,10'h014,8'h43};  //alert-> Tdd 
                12'd1024  :cmd_data={1'b0,10'h017,8'h00};
                default:  cmd_data={1'b0,10'h017,8'h00};
            endcase 
    end
endmodule
